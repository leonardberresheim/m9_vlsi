library ieee;
use ieee.std_logic_1164.all;

entity m9_artan_rom is
    port (i : in std_logic_vector(4 downto 0);
          d : out std_logic_vector(31 downto 0));
end m9_artan_rom;

architecture behaviour of m9_artan_rom is

begin
    with i select d <= 
    "00101101"&"000000000000000000000000" when "00000",
    "00011010"&"100100001010011100110001" when "00001",
    "00001110"&"000010010100011101000000" when "00010",
    "00000111"&"001000000000000100010010" when "00011",
    "00000011"&"100100111000101010100110" when "00100",
    "00000001"&"110010100011011110010100" when "00101",
    "00000000"&"111001010010101000011010" when "00110",
    "00000000"&"011100101001011011010111" when "00111",
    "00000000"&"001110010100101110100101" when "01000",
    "00000000"&"000111001010010111011001" when "01001",
    "00000000"&"000011100101001011101101" when "01010",
    "00000000"&"000001110010100101110110" when "01011",
    "00000000"&"000000111001010010111011" when "01100",
    "00000000"&"000000011100101001011101" when "01101",
    "00000000"&"000000001110010100101110" when "01110",
    "00000000"&"000000000111001010010111" when "01111",
    "00000000"&"000000000011100101001011" when "10000",
    "00000000"&"000000000001110010100101" when "10001",
    "00000000"&"000000000000111001010010" when "10010",
    "00000000"&"000000000000011100101001" when "10011",
    "00000000"&"000000000000001110010100" when "10100",
    "00000000"&"000000000000000111001010" when "10101",
    "00000000"&"000000000000000011100101" when "10110",
    "00000000"&"000000000000000001110010" when "10111",
    "00000000"&"000000000000000000111001" when "11000",
    "00000000"&"000000000000000000011100" when "11001",
    "00000000"&"000000000000000000001110" when "11010",
    "00000000"&"000000000000000000000111" when "11011",
    "00000000"&"000000000000000000000011" when "11100",
    "00000000"&"000000000000000000000001" when "11101",
    "00000000"&"000000000000000000000000" when "11110",
    "00000000"&"000000000000000000000000" when others;

end behaviour;